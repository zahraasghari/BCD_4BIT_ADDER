LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY BCD_4BIT_ADDER IS
PORT(A0,A1,A2,A3,B0,B1,B2,B3:IN STD_LOGIC;
     CIN:IN STD_LOGIC;
	  S0,S1,S2,S3:OUT STD_LOGIC;
       CARRY:OUT STD_LOGIC);
END BCD_4BIT_ADDER;

ARCHITECTURE BCD_4BIT_ADDER_ARCH OF BCD_4BIT_ADDER IS
COMPONENT BITFULLADDER
PORT(A,B,CIN:IN STD_LOGIC;SUM,CARRY:OUT STD_LOGIC);
END COMPONENT;

COMPONENT XOR1
PORT(A,B:IN STD_LOGIC; C:OUT STD_LOGIC);
END COMPONENT;

SIGNAL J0,J1,J2,J3,C1,C2,C3,C4,C5,C6,CR: STD_LOGIC;

BEGIN
STEP11:BITFULLADDER PORT MAP(A0,B0,CIN,J0,C1);
STEP12:BITFULLADDER PORT MAP(A1,B1,C1,J1,C2);
STEP13:BITFULLADDER PORT MAP(A2,B2,C2,J2,C3);
STEP14:BITFULLADDER PORT MAP(A3,B3,C3,J3,C4);

CR<=(((J3 NAND J2)NAND(J3 NAND J1)) NAND ((C4 NAND C4)));
S0<=J0;
STEP15:BITFULLADDER PORT MAP(J1,CR,'0',S1,C5);
STEP16:BITFULLADDER PORT MAP(J2,CR,'0',S2,C6);

STEP21: XOR1 PORT MAP(J3,C6,S3);
CARRY<=CR;


END BCD_4BIT_ADDER_ARCH;