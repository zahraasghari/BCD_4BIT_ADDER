LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY BITFULLADDER IS
PORT(A,B,CIN:IN STD_LOGIC;SUM,CARRY:OUT STD_LOGIC);
END BITFULLADDER;
ARCHITECTURE BITFULLADDER_ARCH OF BITFULLADDER IS
COMPONENT HALF_ADDER
PORT(A,B:IN STD_LOGIC;SUM,CARRY:OUT STD_LOGIC);
END COMPONENT;
SIGNAL Z1,C1,C2: STD_LOGIC;
BEGIN
STEP5:HALF_ADDER PORT MAP(A,B,Z1,C1);
STEP6:HALF_ADDER PORT MAP(CIN,Z1,SUM,C2);
CARRY<=((C1 NAND C1) NAND (C2 NAND C2));
END BITFULLADDER_ARCH;